module helper

